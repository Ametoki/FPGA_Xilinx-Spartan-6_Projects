`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:30:07 06/04/2019 
// Design Name: 
// Module Name:    F20190604 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module F20190604(
    input ext_clk_25m,
    input ext_rst_n,
    output clk_12m5
    );


endmodule
