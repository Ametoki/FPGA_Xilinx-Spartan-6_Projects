`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:28:08 06/09/2019 
// Design Name: 
// Module Name:    SEG_Scan 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module SEG_Scan(
	input           clk,
	input           rst_n,
	output reg[5:0] seg_sel,
	output reg[7:0] seg_data,
	//input[5:0]      seg_en,
	input[7:0]      seg_data_0,
	input[7:0]      seg_data_1,
	input[7:0]      seg_data_2,
	input[7:0]      seg_data_3,
	input[7:0]      seg_data_4,
	input[7:0]      seg_data_5
    );

parameter SCAN_FREQ  = 32'd200;
parameter CLK_FREQ   = 32'd50_000_000;
parameter SCAN_COUNT = CLK_FREQ / (SCAN_FREQ * 6) - 1;

reg[31:0] scan_timer;
reg[3:0]  scan_sel;

always@(posedge clk or negedge rst_n)
begin
	if(!rst_n)
	begin
		scan_timer <= 32'd0;
		scan_sel <= 4'd0;
	end
	else if(scan_timer >= SCAN_COUNT)
	begin
		scan_timer <= 32'd0;
		if(scan_sel == 4'd5)
			scan_sel <= 4'd0;
		else
			scan_sel <= scan_sel + 4'd1;
	end
	else
		begin
			scan_timer <= scan_timer + 32'd1;
		end
end
always@(posedge clk or negedge rst_n)
begin
	if(!rst_n)
	begin
		seg_sel <= 6'b111_111;
		seg_data <= 8'hff;
	end
	else
	begin
		case(scan_sel)
			4'd0:
			begin
				seg_sel  <= 6'b11_1110;
				seg_data <= seg_data_0;
			end
			4'd1:
			begin
				seg_sel  <= 6'b11_1101;
				seg_data <= seg_data_1;
			end
			4'd2:
			begin
				seg_sel  <= 6'b11_1011;
				seg_data <= seg_data_2;
			end
			4'd3:
			begin
				seg_sel  <= 6'b11_0111;
				seg_data <= seg_data_3;
			end
			4'd4:
			begin
				seg_sel  <= 6'b10_1111;
				seg_data <= seg_data_4;
			end
			4'd5:
			begin
				seg_sel  <= 6'b01_1111;
				seg_data <= seg_data_5;
			end
			default:
			begin
				seg_sel  <= 6'b11_1111;
				seg_data <= 8'hff;
			end
		endcase
	end
end

endmodule
